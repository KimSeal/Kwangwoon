module _XOR(A,B,Y);//XOR function
	input A,B;
	output Y;
	assign Y = A ^ B;//^ equals (+)
endmodule
