library verilog;
use verilog.vl_types.all;
entity tb_XOR is
end tb_XOR;
